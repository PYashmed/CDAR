//˫ɫ�����ۺ�����ģ��
//����mode��00xxΪcat��xx֡����������00-11 01xx��dog  10xx��mouse






module dotmatric (
    input clk1khz,output [7:0]row,colr,colg,input [3:0]mode,input rst,off
);
    wire [7:0]cat,dog,mouse;
    wire [2:0]cnt;
    cnt8 u1(
        .clk(clk1khz),
        .cnt(cnt)
    );
    bicolor_dot_matrix u2(
        .cnt(cnt),
        .row(row),
        .r(colr),
        .g(colg),
        .cat(cat),
        .dog(dog),
        .mouse(mouse),
        .off(off)
    );

    changemode u3(
        .mode(mode),
        .clk1hz(clk1hz),
        .cat(cat),
        .dog(dog),
        .mouse(mouse),
        .rst(rst)
    );
    divide #(.wide(10),.n(500)) u4(
        .clk(clk1khz),
        .clkout(clk1hz)
    );
endmodule
//��ɨ�����ʱ�ӣ�����ģ�飩
module cnt8 (
    input clk,output reg [2:0]cnt
);
always @(posedge clk) begin
    if(cnt==3'b111)
        cnt=3'b000;
    else
        cnt=cnt+1'b1;
end
endmodule



//��������ģ��(��ɨ����ʾ)
module bicolor_dot_matrix (
    output reg [7:0]r,g,row,input [2:0]cnt,input [7:0]cat,dog,mouse,input off
);
//��ʾģ�飨��ɨ����ʾ��
always @(cnt) begin
    if(off)begin
        row<=8'b11111111;
    end
    else begin
        case(cnt)
            3'b000:begin row<=8'b11111110;r<=cat; g<=8'b0; end
            3'b001:begin row<=8'b11111101;r<=cat; g<=8'b0; end
            3'b010:begin row<=8'b11111011;r<=8'b0; g<=8'b0; end
            3'b011:begin row<=8'b11110111;r<=8'b0; g<=dog; end
            3'b100:begin row<=8'b11101111;r<=8'b0; g<=dog; end
            3'b101:begin row<=8'b11011111;r<=8'b0;g<=8'b0; end
            3'b110:begin row<=8'b10111111;r<=mouse;g<=mouse; end
            3'b111:begin row<=8'b01111111;r<=mouse;g<=mouse; end
            default:row<=8'b11111111;
        endcase
    end
end
endmodule


module changemode (
    input [3:0]mode,output reg [7:0]cat,dog,mouse,input clk1hz,rst
);

initial begin
    cat=8'b11000000;
    dog=8'b11000000;
    mouse=8'b11000000;
end
//����ÿ֡
always @(posedge clk1hz or posedge rst) begin
    if(rst)begin
        cat<=8'b11000000;
        dog<=8'b11000000;
        mouse<=8'b11000000;
    end
    else begin

        case(mode)//ǰ��λ��00��cat 01��dog 10��mouse������λ��00��0֡��ԭλ�ã�01��1֡ 10��2֡ 11��3֡
            4'b0000:begin cat<=8'b11000000; dog<=dog; mouse<=mouse; end
            4'b0001:begin cat<=8'b00110000; dog<=dog; mouse<=mouse; end
            4'b0010:begin cat<=8'b00001100; dog<=dog; mouse<=mouse; end
            4'b0011:begin cat<=8'b00000011; dog<=dog; mouse<=mouse; end
            4'b0100:begin cat<=cat; dog<=8'b11000000; mouse<=mouse; end
            4'b0101:begin cat<=cat; dog<=8'b00110000; mouse<=mouse; end
            4'b0110:begin cat<=cat; dog<=8'b00001100; mouse<=mouse; end
            4'b0111:begin cat<=cat; dog<=8'b00000011; mouse<=mouse; end
            4'b1000:begin cat<=cat; dog<=dog; mouse<=8'b11000000; end
            4'b1001:begin cat<=cat; dog<=dog; mouse<=8'b00110000; end
            4'b1010:begin cat<=cat; dog<=dog; mouse<=8'b00001100; end
            4'b1011:begin cat<=cat; dog<=dog; mouse<=8'b00000011; end
            default:begin cat<=cat; dog<=dog; mouse<=mouse; end
        endcase
    end
end

endmodule


module divide (input clk,output clkout);
	parameter	wide = 3;
	parameter	n = 5;
 
	reg [wide-1:0]	cntp,cntn;
	reg clkp,clkn;
	//�����ش���ʱ�������Ŀ���
always @(posedge clk)
	begin
		if (cntp==(n-1))
			cntp<=0;
		else cntp<=cntp+1;//ģn�ļ�����
	end

	//�����ش����ķ�Ƶʱ�����,���nΪ�����õ���ʱ��ռ�ձȲ���50%�����nΪż���õ���ʱ��ռ�ձ�Ϊ50%
always @(posedge clk)
	begin
		if (cntp<(n>>1))//����2ȥ������
			clkp<=0;
		else 
			clkp<=1;//�õ��ķ�Ƶʱ�������ڱȸ����ڶ�һ��clkʱ��
	end

	//�½��ش���ʱ�������Ŀ���
always @(negedge clk)
	begin
		if (cntn==(n-1))
			cntn<=0;
		else cntn<=cntn+1;
	end

	//�½��ش����ķ�Ƶʱ���������clkp�����ʱ��
always @(negedge clk)
	begin
		if (cntn<(n>>1))  
			clkn<=0;
		else 
			clkn<=1;//�õ��ķ�Ƶʱ�������ڱȸ����ڶ�һ��clkʱ��
	end

    assign clkout = (n==1)?clk:(n[0])?(clkp&clkn):clkp;//�����жϱ��ʽ
                                                          //��n=1ʱ��ֱ�����clk
                                                          //��nΪż��Ҳ����n�����λΪ0��n��0��=0�����clkp
                                                          //��nΪ����Ҳ����n���λΪ1��n��0��=1�����clkp&clkn�������ڶ�����������
endmodule