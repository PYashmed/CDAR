module game (
    
);
    


    
endmodule